LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY UART IS
	PORT(
		
	);
END ENTITY;

ARCHITECTURE behavior OF UART IS
BEGIN
	
END ARCHITECTURE;