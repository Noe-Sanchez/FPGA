library IEEE;
use IEEE.std_logic_1164.all;

entity equipo4_fsm_3_1 is
    port(
        clk, rst :   in      std_logic;
    	ab       :   in      std_logic_vector(1 downto 0);
    	z        :   out     std_logic
    );
end entity;

architecture behaviour of equipo4_fsm_3_1 is
    signal c_state  :   std_logic_vector(2 downto 0) := "000";
    signal a, b   :     std_logic;
begin
    process(clk)
        begin
            a <= ab(1);
            b <= ab(0);
            if clk = '1' then
                if rst = '1' then
                    z <= '0';
                    c_state <= "000";
                elsif c_state = "000" then
                        z <= '0';
                        if (a='1') and (b='1') then
                            c_state <= "001";
                        end if;   
                elsif c_state = "001" then
                    z <= '0';
                    if a='0' and b='1' then
                        c_state <= "010";
                    elsif a='1' and b='0' then
                        c_state <= "000";
                    end if;
                elsif c_state = "010" then
                    z <= '1';
                    if a='1' or b='1' then
                        c_state <= "011";
                    end if;
                elsif c_state = "100" then
                    z <= '0';
                    c_state <= "000";
                else
                    c_state <= "000";
                end if;
            end if;
        end process;
end architecture;


  
